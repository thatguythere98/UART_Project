`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:
// Design Name:
// Module Name:
// Project Name:
// Target Devices:
// Tool Versions:
// Description: Testbench, not up to date.
//
// Dependencies: 
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module tb_Tx;

  // Inputs
  reg        clk;  // Clock signal
  reg        rst;  // Active-low reset signal
  reg  [7:0] din;  // Data input
  reg        tx_start;  // Transmission start signal

  // Outputs
  wire       tx;  // UART transmit output
  wire       tx_done;  // Transmission done signal
  wire       sample_clk;  // 16x Baud rate clock, generated by BaudGenerator


  // Instantiate the Unit Under Test (UUT)
  Tx Dut (
       .clk(clk),
       .rst(rst),
       .din(din),
       .tx_start(tx_start),
       .sample_tick(sample_clk),
       .tx(tx),
       .tx_done(tx_done)
     );
  // Instantiate the BaudGenerator module
  BaudGenerator baud_gen (
                  .rst(rst),
                  .clk(clk),
                  .sel(3'b000),       // Set to 9600 baud for this example
                  .baud16x_out(sample_clk)  // Connect baud16x_out to sample_clk
                );

  initial
  begin
    clk = 0;
    forever
      #41.660 clk = ~clk;  // 7.3728 MHz clock
  end

  initial
  begin
    // Initialize Inputs
    clk      = 0;  // Initial clock state
    rst      = 1;  // Assert reset
    din      = 8'b0;  // Clear data input
    tx_start = 0;  // Clear start signal

    // Apply reset
    #20;
    rst      = 0;  // Deassert reset

    // Test case: Transmit 0x6A, FF
    din      = 8'b00001111;  // Set data to 0x45
    tx_start = 1;  // Assert start signal
    #600;
    tx_start = 0;  // Deassert start signal

    // Wait for transmission to complete
    wait (tx_done);  // Wait until transmission is done
    #40;  // Wait some time before next test

    // Test case: Transmit 0x96
    din      = 8'b11110000;  // Set data to 0x18
    tx_start = 1;  // Assert start signal
    #600;
    tx_start = 0;  // Deassert start signal

    // Wait for transmission to complete
    wait (tx_done);  // Wait until transmission is done
    #40;  // Wait some time before ending simulation

    // End simulation
    $stop;  // Stop the simulation
  end
endmodule
