`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:
// Design Name:
// Module Name:
// Project Name:
// Target Devices:
// Tool Versions:
// Description: Testbench, not up to date.
//
// Dependencies: 
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module tb_Rx;

  // Testbench signals
  reg clk;           // System clock (for BaudGenerator)
  reg rst;
  reg rx;
  wire sample_clk;   // 16x Baud rate clock, generated by BaudGenerator
  wire [7:0] dout;
  wire rx_done;

  // Instantiate the Rx module
  Rx Dut (
       .clk(clk),
       .rst(rst),
       .rx(rx),
       .sample_tick(sample_clk),  // Connect baud16x_out to sample_tick
       .dout(dout),
       .rx_done(rx_done)
     );

  // Instantiate the BaudGenerator module
  BaudGenerator baud_gen (
                  .rst(rst),
                  .clk(clk),
                  .sel(3'b000),       // Set to 9600 baud for this example
                  .baud16x_out(sample_clk)  // Connect baud16x_out to sample_clk
                );


  initial
  begin
    clk = 0;
    forever
     #67.815 clk = ~clk;  // 7.3728 MHz clock
  end

  // Test stimulus
  initial
  begin
    // Initialize signals
    rst = 0;
    rx = 1;

    // Apply reset
    #100;
    rst = 1;
    #100;
    rst = 0;
    #100;

    // Send a byte: 0xA5 (0b10100101)
    send_byte(8'b10100101); //0xA5
    send_byte(8'b11111111); //xFF
    send_byte(8'b01010101); //0x55

    // Wait for reception to complete
    #200000;
    if (dout == 8'b10100101 && rx_done)
    begin
      $display("Test Passed: Received byte 0xA5 correctly.");
    end
    else
    begin
      $display("Test Failed: Incorrect byte received.");
    end

    // End of simulation
    $finish;
  end

  // Task to send a byte over UART
  task send_byte(input [7:0] byteData);
    integer i;
    begin
      // Send start bit
      rx = 0;
      #(104167);  // Wait one bit period (baud rate clock)

      // Send data bits (LSB first)
      for (i = 0; i < 8; i = i + 1)
      begin
        rx = byteData[i];
        #(104167);  // Wait one bit period
      end

      // Send stop bit
      rx = 1;
      #(104167);  // Wait one bit period

      // Ensure idle line
      #(104167);
    end
  endtask

endmodule